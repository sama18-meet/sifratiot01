// Full Adder/Subtractor test bench template
module fas_test;

// Put your code here
// ------------------


// End of your code

endmodule
