// 4->1 multiplexer test bench template
module mux4_test;

// Put your code here
// ------------------


// End of your code

endmodule
